Eight_Bit_Divider_inst : Eight_Bit_Divider PORT MAP (
		aclr	 => aclr_sig,
		clken	 => clken_sig,
		clock	 => clock_sig,
		denom	 => denom_sig,
		numer	 => numer_sig,
		quotient	 => quotient_sig,
		remain	 => remain_sig
	);
