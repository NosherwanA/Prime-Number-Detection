library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity MRT is
    port(

    );
end entity;

architecture internal of MRT is



    begin



end architecture;